//: version "1.8.7"

module HA(C, S, B, A);
//: interface  /sz:(72, 76) /bd:[ Ti0>B(58/72) Ti1>A(19/72) Lo0<C(37/76) Bo0<S(28/72) ]
input B;    //: /sn:0 {0}(122,340)(208,340){1}
//: {2}(212,340)(257,340)(257,326)(265,326){3}
//: {4}(210,342)(210,371)(265,371){5}
input A;    //: /sn:0 {0}(122,321)(225,321){1}
//: {2}(229,321)(265,321){3}
//: {4}(227,323)(227,366)(265,366){5}
output C;    //: /sn:0 /dp:1 {0}(286,369)(380,369){1}
output S;    //: /sn:0 /dp:1 {0}(286,324)(375,324){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(276,324) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  //: output g3 (C) @(377,369) /sn:0 /w:[ 1 ]
  //: output g2 (S) @(372,324) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(120,340) /sn:0 /w:[ 0 ]
  //: joint g6 (B) @(210, 340) /w:[ 2 -1 1 4 ]
  //: joint g7 (A) @(227, 321) /w:[ 2 -1 1 4 ]
  and g5 (.I0(A), .I1(B), .Z(C));   //: @(276,369) /sn:0 /delay:" 3" /w:[ 5 5 0 ]
  //: input g0 (A) @(120,321) /sn:0 /w:[ 0 ]

endmodule

module RCA(S, B, A);
//: interface  /sz:(113, 97) /bd:[ Ti0>A[3:0](38/113) Ti1>B[3:0](75/113) Bo0<S[7:0](53/113) ]
input [3:0] B;    //: /sn:0 /dp:9 {0}(659,463)(659,447){1}
//: {2}(659,446)(659,247){3}
//: {4}(659,246)(659,83){5}
//: {6}(659,82)(659,36){7}
//: {8}(659,35)(659,9){9}
input [3:0] A;    //: /sn:0 {0}(-20,26)(6,26)(6,12){1}
//: {2}(6,11)(6,3){3}
//: {4}(6,2)(6,-6){5}
//: {6}(6,-7)(6,-14){7}
//: {8}(6,-15)(6,-21){9}
output [7:0] S;    //: /sn:0 /dp:1 {0}(625,675)(674,675)(674,677)(683,677){1}
wire w6;    //: /sn:0 {0}(567,72)(567,640)(619,640){1}
wire w13;    //: /sn:0 /dp:1 {0}(-39,382)(-117,382)(-117,504){1}
wire w7;    //: /sn:0 {0}(10,3)(106,3){1}
//: {2}(110,3)(155,3){3}
//: {4}(159,3)(231,3){5}
//: {6}(235,3)(319,3)(319,48){7}
//: {8}(233,5)(233,104){9}
//: {10}(157,5)(157,277){11}
//: {12}(108,5)(108,135)(52,135)(52,437)(30,437)(30,458){13}
wire w50;    //: /sn:0 {0}(221,227)(221,324)(196,324)(196,339){1}
wire w34;    //: /sn:0 {0}(84,121)(84,149){1}
wire w4;    //: /sn:0 {0}(215,416)(215,494)(221,494)(221,504){1}
wire w39;    //: /sn:0 {0}(236,125)(236,150){1}
wire w56;    //: /sn:0 {0}(484,126)(484,151){1}
wire w3;    //: /sn:0 {0}(178,380)(143,380){1}
wire w0;    //: /sn:0 {0}(10,12)(33,12){1}
//: {2}(37,12)(59,12){3}
//: {4}(63,12)(79,12){5}
//: {6}(83,12)(199,12)(199,48){7}
//: {8}(81,14)(81,100){9}
//: {10}(61,14)(61,118)(-86,118)(-86,462){11}
//: {12}(35,14)(35,276){13}
wire w22;    //: /sn:0 {0}(10,-6)(173,-6){1}
//: {2}(177,-6)(268,-6){3}
//: {4}(272,-6)(350,-6){5}
//: {6}(354,-6)(441,-6)(441,49){7}
//: {8}(352,-4)(352,105){9}
//: {10}(270,-4)(270,282){11}
//: {12}(175,-4)(175,341)(161,341)(161,433)(144,433)(144,459){13}
wire w60;    //: /sn:0 {0}(147,480)(147,502){1}
wire w20;    //: /sn:0 {0}(38,297)(38,316)(13,316)(13,341){1}
wire w29;    //: /sn:0 {0}(132,579)(132,680)(619,680){1}
wire w42;    //: /sn:0 {0}(298,379)(250,379){1}
wire w12;    //: /sn:0 {0}(109,227)(109,315)(89,315)(89,340){1}
wire w19;    //: /sn:0 {0}(-98,581)(-98,700)(619,700){1}
wire w18;    //: /sn:0 /dp:1 {0}(-135,545)(-145,545)(-145,710)(619,710){1}
wire w66;    //: /sn:0 {0}(-83,483)(-83,504){1}
wire w23;    //: /sn:0 {0}(-19,544)(-63,544){1}
wire w63;    //: /sn:0 {0}(33,479)(33,503){1}
wire w54;    //: /sn:0 {0}(303,190)(256,190){1}
wire w21;    //: /sn:0 {0}(202,69)(202,150){1}
wire w24;    //: /sn:0 {0}(18,580)(18,690)(619,690){1}
wire w31;    //: /sn:0 {0}(388,300)(388,320)(357,320)(357,341){1}
wire w32;    //: /sn:0 {0}(201,542)(167,542){1}
wire w53;    //: /sn:0 {0}(654,83)(488,83){1}
//: {2}(484,83)(359,83){3}
//: {4}(355,83)(240,83){5}
//: {6}(236,83)(86,83)(86,100){7}
//: {8}(238,85)(238,104){9}
//: {10}(357,85)(357,105){11}
//: {12}(486,85)(486,105){13}
wire w8;    //: /sn:0 {0}(71,381)(33,381){1}
wire w52;    //: /sn:0 /dp:1 {0}(-81,462)(-81,447)(33,447){1}
//: {2}(37,447)(147,447){3}
//: {4}(151,447)(260,447){5}
//: {6}(264,447)(654,447){7}
//: {8}(262,449)(262,463){9}
//: {10}(149,449)(149,459){11}
//: {12}(35,449)(35,458){13}
wire w27;    //: /sn:0 {0}(322,69)(322,139)(321,139)(321,149){1}
wire w44;    //: /sn:0 {0}(425,189)(375,189){1}
wire w17;    //: /sn:0 {0}(40,276)(40,247)(160,247){1}
//: {2}(164,247)(273,247){3}
//: {4}(277,247)(388,247){5}
//: {6}(392,247)(654,247){7}
//: {8}(390,249)(390,279){9}
//: {10}(275,249)(275,282){11}
//: {12}(162,249)(162,277){13}
wire w35;    //: /sn:0 {0}(444,70)(444,141)(445,141)(445,151){1}
wire w33;    //: /sn:0 {0}(246,582)(246,670)(619,670){1}
wire w28;    //: /sn:0 {0}(95,543)(53,543){1}
wire w45;    //: /sn:0 {0}(470,229)(470,650)(619,650){1}
wire w49;    //: /sn:0 {0}(184,191)(138,191){1}
wire w14;    //: /sn:0 {0}(-2,418)(-2,493)(-1,493)(-1,503){1}
wire w2;    //: /sn:0 {0}(654,36)(571,36){1}
//: {2}(567,36)(448,36){3}
//: {4}(444,36)(326,36){5}
//: {6}(322,36)(204,36)(204,48){7}
//: {8}(324,38)(324,48){9}
//: {10}(446,38)(446,49){11}
//: {12}(569,38)(569,51){13}
wire w11;    //: /sn:0 {0}(64,187)(-21,187)(-21,341){1}
wire w48;    //: /sn:0 {0}(355,126)(355,149){1}
wire w47;    //: /sn:0 {0}(160,298)(160,314)(123,314)(123,340){1}
wire w55;    //: /sn:0 {0}(340,226)(340,320)(318,320)(318,341){1}
wire w38;    //: /sn:0 {0}(273,303)(273,323)(230,323)(230,339){1}
wire w43;    //: /sn:0 {0}(343,419)(343,660)(619,660){1}
wire w9;    //: /sn:0 {0}(108,417)(108,492)(113,492)(113,502){1}
wire w26;    //: /sn:0 {0}(10,-14)(285,-14){1}
//: {2}(289,-14)(383,-14){3}
//: {4}(387,-14)(479,-14){5}
//: {6}(483,-14)(564,-14)(564,51){7}
//: {8}(481,-12)(481,105){9}
//: {10}(385,-12)(385,279){11}
//: {12}(287,-12)(287,431)(257,431)(257,463){13}
wire w57;    //: /sn:0 {0}(260,484)(260,504){1}
//: enddecls

  FA g8 (.A(w9), .B(w60), .Cin(w32), .Cout(w28), .S(w29));   //: @(96, 503) /sz:(70, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  FA g4 (.A(w12), .B(w47), .Cin(w3), .Cout(w8), .S(w9));   //: @(72, 341) /sz:(70, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  and g44 (.I0(w7), .I1(w52), .Z(w63));   //: @(33,469) /sn:0 /R:3 /delay:" 3" /w:[ 13 13 0 ]
  and g16 (.I0(w0), .I1(w2), .Z(w21));   //: @(202,59) /sn:0 /R:3 /delay:" 3" /w:[ 7 7 0 ]
  FA g3 (.A(w50), .B(w38), .Cin(w42), .Cout(w3), .S(w4));   //: @(179, 340) /sz:(70, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  and g47 (.I0(w0), .I1(w17), .Z(w20));   //: @(38,287) /sn:0 /R:3 /delay:" 3" /w:[ 13 0 0 ]
  and g17 (.I0(w7), .I1(w2), .Z(w27));   //: @(322,59) /sn:0 /R:3 /delay:" 3" /w:[ 7 9 0 ]
  //: joint g26 (w2) @(569, 36) /w:[ 1 -1 2 12 ]
  //: output g2 (S) @(680,677) /sn:0 /w:[ 1 ]
  tran g23(.Z(w2), .I(B[0]));   //: @(657,36) /sn:0 /R:2 /w:[ 0 7 8 ] /ss:0
  and g30 (.I0(w26), .I1(w53), .Z(w56));   //: @(484,116) /sn:0 /R:3 /delay:" 3" /w:[ 9 13 0 ]
  //: input g1 (B) @(659,7) /sn:0 /R:3 /w:[ 9 ]
  //: joint g24 (w2) @(324, 36) /w:[ 5 -1 6 8 ]
  and g39 (.I0(w26), .I1(w17), .Z(w31));   //: @(388,290) /sn:0 /R:3 /delay:" 3" /w:[ 11 9 0 ]
  and g29 (.I0(w22), .I1(w53), .Z(w48));   //: @(355,116) /sn:0 /R:3 /delay:" 3" /w:[ 9 11 0 ]
  //: joint g60 (w22) @(175, -6) /w:[ 2 -1 1 12 ]
  //: joint g51 (w17) @(162, 247) /w:[ 2 -1 1 12 ]
  and g18 (.I0(w22), .I1(w2), .Z(w35));   //: @(444,60) /sn:0 /R:3 /delay:" 3" /w:[ 7 11 0 ]
  HA g10 (.A(w34), .B(w49), .C(w11), .S(w12));   //: @(65, 150) /sz:(72, 76) /sn:0 /p:[ Ti0>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g25 (w2) @(446, 36) /w:[ 3 -1 4 10 ]
  //: joint g49 (w17) @(390, 247) /w:[ 6 -1 5 8 ]
  FA g6 (.A(w13), .B(w66), .Cin(w23), .Cout(w18), .S(w19));   //: @(-134, 505) /sz:(70, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g50 (w17) @(275, 247) /w:[ 4 -1 3 10 ]
  HA g9 (.A(w4), .B(w57), .C(w32), .S(w33));   //: @(202, 505) /sz:(72, 76) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<0 ]
  FA g7 (.A(w14), .B(w63), .Cin(w28), .Cout(w23), .S(w24));   //: @(-18, 504) /sz:(70, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g35 (w0) @(81, 12) /w:[ 6 -1 5 8 ]
  //: joint g56 (w52) @(35, 447) /w:[ 2 -1 1 12 ]
  //: joint g58 (w52) @(262, 447) /w:[ 6 -1 5 8 ]
  tran g31(.Z(w53), .I(B[1]));   //: @(657,83) /sn:0 /R:2 /w:[ 0 5 6 ] /ss:0
  tran g22(.Z(w0), .I(A[3]));   //: @(4,12) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:1
  //: joint g59 (w26) @(287, -14) /w:[ 2 -1 1 12 ]
  //: joint g33 (w53) @(357, 83) /w:[ 3 -1 4 10 ]
  //: joint g36 (w7) @(233, 3) /w:[ 6 -1 5 8 ]
  and g41 (.I0(w7), .I1(w17), .Z(w47));   //: @(160,288) /sn:0 /R:3 /delay:" 3" /w:[ 11 13 0 ]
  and g45 (.I0(w0), .I1(w52), .Z(w66));   //: @(-83,473) /sn:0 /R:3 /delay:" 3" /w:[ 11 0 0 ]
  //: joint g54 (w7) @(157, 3) /w:[ 4 -1 3 10 ]
  and g40 (.I0(w22), .I1(w17), .Z(w38));   //: @(273,293) /sn:0 /R:3 /delay:" 3" /w:[ 11 11 0 ]
  and g42 (.I0(w26), .I1(w52), .Z(w57));   //: @(260,474) /sn:0 /R:3 /delay:" 3" /w:[ 13 9 0 ]
  //: joint g52 (w26) @(385, -14) /w:[ 4 -1 3 10 ]
  HA g12 (.A(w35), .B(w56), .C(w44), .S(w45));   //: @(426, 152) /sz:(72, 76) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<0 ]
  and g28 (.I0(w7), .I1(w53), .Z(w39));   //: @(236,115) /sn:0 /R:3 /delay:" 3" /w:[ 9 9 0 ]
  //: joint g34 (w53) @(486, 83) /w:[ 1 -1 2 12 ]
  tran g46(.Z(w17), .I(B[2]));   //: @(657,247) /sn:0 /R:2 /w:[ 7 3 4 ] /ss:0
  //: joint g57 (w52) @(149, 447) /w:[ 4 -1 3 10 ]
  FA g14 (.A(w27), .B(w48), .Cin(w44), .Cout(w54), .S(w55));   //: @(304, 150) /sz:(70, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  FA g5 (.A(w11), .B(w20), .Cin(w8), .Cout(w13), .S(w14));   //: @(-38, 342) /sz:(70, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  HA g11 (.A(w55), .B(w31), .C(w42), .S(w43));   //: @(299, 342) /sz:(72, 76) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<0 ]
  tran g19(.Z(w26), .I(A[0]));   //: @(4,-14) /sn:0 /R:2 /w:[ 0 7 8 ] /ss:1
  tran g21(.Z(w7), .I(A[2]));   //: @(4,3) /sn:0 /R:2 /w:[ 0 3 4 ] /ss:1
  //: joint g61 (w7) @(108, 3) /w:[ 2 -1 1 12 ]
  //: joint g32 (w53) @(238, 83) /w:[ 5 -1 6 8 ]
  tran g20(.Z(w22), .I(A[1]));   //: @(4,-6) /sn:0 /R:2 /w:[ 0 5 6 ] /ss:1
  concat g63 (.I0(w6), .I1(w45), .I2(w43), .I3(w33), .I4(w29), .I5(w24), .I6(w19), .I7(w18), .Z(S));   //: @(624,675) /sn:0 /w:[ 1 1 1 1 1 1 1 1 0 ] /dr:1
  and g15 (.I0(w26), .I1(w2), .Z(w6));   //: @(567,62) /sn:0 /R:3 /delay:" 3" /w:[ 7 13 0 ]
  //: input g0 (A) @(-22,26) /sn:0 /w:[ 0 ]
  //: joint g38 (w26) @(481, -14) /w:[ 6 -1 5 8 ]
  and g43 (.I0(w22), .I1(w52), .Z(w60));   //: @(147,470) /sn:0 /R:3 /delay:" 3" /w:[ 13 11 0 ]
  and g27 (.I0(w0), .I1(w53), .Z(w34));   //: @(84,111) /sn:0 /R:3 /delay:" 3" /w:[ 9 7 0 ]
  tran g48(.Z(w52), .I(B[3]));   //: @(657,447) /sn:0 /R:2 /w:[ 7 1 2 ] /ss:0
  //: joint g37 (w22) @(352, -6) /w:[ 6 -1 5 8 ]
  //: joint g62 (w0) @(61, 12) /w:[ 4 -1 3 10 ]
  //: joint g55 (w0) @(35, 12) /w:[ 2 -1 1 12 ]
  FA g13 (.A(w21), .B(w39), .Cin(w54), .Cout(w49), .S(w50));   //: @(185, 151) /sz:(70, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g53 (w22) @(270, -6) /w:[ 4 -1 3 10 ]

endmodule

module FA(Cout, S, Cin, B, A);
//: interface  /sz:(70, 75) /bd:[ Ti0>B(51/70) Ti1>A(17/70) Ri0>Cin(39/75) Lo0<Cout(40/75) Bo0<S(34/70) ]
input B;    //: /sn:0 {0}(125,198)(216,198){1}
input A;    //: /sn:0 {0}(125,181)(216,181){1}
input Cin;    //: /sn:0 {0}(132,107)(277,107){1}
output Cout;    //: /sn:0 /dp:1 {0}(392,153)(419,153){1}
output S;    //: /sn:0 {0}(299,98)(299,67)(317,67){1}
wire w1;    //: /sn:0 {0}(239,175)(239,155)(371,155){1}
wire w8;    //: /sn:0 {0}(259,199)(269,199)(269,121)(277,121){1}
wire w5;    //: /sn:0 {0}(319,114)(361,114)(361,150)(371,150){1}
//: enddecls

  //: output g4 (Cout) @(416,153) /sn:0 /w:[ 1 ]
  //: output g3 (S) @(314,67) /sn:0 /w:[ 1 ]
  //: input g2 (Cin) @(130,107) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(123,198) /sn:0 /w:[ 0 ]
  HA g6 (.B(w8), .A(Cin), .S(S), .C(w5));   //: @(278, 99) /sz:(40, 40) /sn:0 /p:[ Li0>1 Li1>1 To0<0 Ro0<0 ]
  or g9 (.I0(w5), .I1(w1), .Z(Cout));   //: @(382,153) /sn:0 /delay:" 3" /w:[ 1 1 0 ]
  HA g5 (.B(B), .A(A), .C(w1), .S(w8));   //: @(217, 176) /sz:(41, 40) /sn:0 /p:[ Li0>1 Li1>1 To0<0 Ro0<0 ]
  //: input g0 (A) @(123,181) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire [3:0] w4;    //: /sn:0 /dp:1 {0}(358,91)(358,151)(301,151)(301,161){1}
wire [3:0] w3;    //: /sn:0 /dp:1 {0}(207,93)(207,151)(264,151)(264,161){1}
wire [7:0] w2;    //: /sn:0 {0}(279,260)(279,284){1}
//: {2}(281,286)(355,286)(355,306){3}
//: {4}(277,286)(210,286)(210,320)(227,333)(185,333){5}
//: {6}(279,288)(279,332){7}
//: enddecls

  led g4 (.I(w2));   //: @(355,313) /sn:0 /R:2 /w:[ 3 ] /type:1
  led g3 (.I(w2));   //: @(279,339) /sn:0 /R:2 /w:[ 7 ] /type:3
  //: dip g2 (w4) @(358,81) /sn:0 /w:[ 0 ] /st:15
  //: dip g1 (w3) @(207,83) /sn:0 /w:[ 0 ] /st:1
  led g6 (.I(w2));   //: @(178,333) /sn:0 /R:1 /w:[ 5 ] /type:2
  //: joint g5 (w2) @(279, 286) /w:[ 2 1 4 6 ]
  RCA g0 (.B(w4), .A(w3), .S(w2));   //: @(226, 162) /sz:(113, 97) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 ]

endmodule
