//: version "1.8.7"

module FA2(Cout, S, Cin, B, A);
//: interface  /sz:(137, 126) /bd:[ Li0>Cin(101/126) Li1>B(66/126) Li2>A(30/126) To0<Cout(72/137) Ro0<S(64/126) ]
input B;    //: /sn:0 {0}(144,181)(144,255){1}
//: {2}(146,257)(218,257){3}
//: {4}(144,259)(144,377){5}
//: {6}(146,379)(159,379)(159,376)(218,376){7}
//: {8}(144,381)(144,415)(218,415){9}
input A;    //: /sn:0 {0}(113,181)(113,239){1}
//: {2}(115,241)(208,241)(208,252)(218,252){3}
//: {4}(113,243)(113,312){5}
//: {6}(115,314)(126,314)(126,323)(219,323){7}
//: {8}(113,316)(113,371)(218,371){9}
input Cin;    //: /sn:0 {0}(173,180)(173,270){1}
//: {2}(175,272)(341,272){3}
//: {4}(173,274)(173,326){5}
//: {6}(175,328)(219,328){7}
//: {8}(173,330)(173,420)(218,420){9}
output Cout;    //: /sn:0 {0}(392,381)(455,381){1}
output S;    //: /sn:0 {0}(362,270)(451,270){1}
wire w8;    //: /sn:0 {0}(240,326)(280,326)(280,337)(325,337){1}
wire w17;    //: /sn:0 {0}(346,340)(361,340)(361,378)(371,378){1}
wire w14;    //: /sn:0 {0}(239,418)(361,418)(361,383)(371,383){1}
wire w2;    //: /sn:0 {0}(239,255)(331,255)(331,267)(341,267){1}
wire w11;    //: /sn:0 {0}(239,374)(283,374)(283,342)(325,342){1}
//: enddecls

  xor g4 (.I0(w2), .I1(Cin), .Z(S));   //: @(352,270) /sn:0 /delay:" 5" /w:[ 1 3 0 ]
  or g8 (.I0(w8), .I1(w11), .Z(w17));   //: @(336,340) /sn:0 /delay:" 4" /w:[ 1 1 0 ]
  xor g3 (.I0(A), .I1(B), .Z(w2));   //: @(229,255) /sn:0 /delay:" 5" /w:[ 3 3 0 ]
  //: output g16 (Cout) @(452,381) /sn:0 /w:[ 1 ]
  //: output g17 (S) @(448,270) /sn:0 /w:[ 1 ]
  //: input g2 (Cin) @(173,178) /sn:0 /R:3 /w:[ 0 ]
  //: input g1 (B) @(144,179) /sn:0 /R:3 /w:[ 0 ]
  //: joint g10 (B) @(144, 379) /w:[ 6 5 -1 8 ]
  and g6 (.I0(A), .I1(B), .Z(w11));   //: @(229,374) /sn:0 /delay:" 4" /w:[ 9 7 0 ]
  and g7 (.I0(B), .I1(Cin), .Z(w14));   //: @(229,418) /sn:0 /delay:" 4" /w:[ 9 9 0 ]
  or g9 (.I0(w17), .I1(w14), .Z(Cout));   //: @(382,381) /sn:0 /delay:" 4" /w:[ 1 1 0 ]
  //: joint g12 (A) @(113, 314) /w:[ 6 5 -1 8 ]
  and g5 (.I0(A), .I1(Cin), .Z(w8));   //: @(230,326) /sn:0 /delay:" 4" /w:[ 7 7 0 ]
  //: joint g11 (Cin) @(173, 328) /w:[ 6 5 -1 8 ]
  //: joint g14 (B) @(144, 257) /w:[ 2 1 -1 4 ]
  //: input g0 (A) @(113,179) /sn:0 /R:3 /w:[ 0 ]
  //: joint g15 (Cin) @(173, 272) /w:[ 2 1 -1 4 ]
  //: joint g13 (A) @(113, 241) /w:[ 2 1 -1 4 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(298,184)(328,184){1}
wire w7;    //: /sn:0 {0}(299,219)(328,219){1}
wire w4;    //: /sn:0 {0}(467,182)(501,182){1}
wire w3;    //: /sn:0 {0}(401,117)(401,98){1}
wire w5;    //: /sn:0 {0}(298,148)(328,148){1}
//: enddecls

  led g4 (.I(w3));   //: @(401,91) /sn:0 /w:[ 1 ] /type:0
  //: switch g3 (w7) @(282,219) /sn:0 /w:[ 0 ] /st:0
  //: switch g2 (w6) @(281,184) /sn:0 /w:[ 0 ] /st:0
  //: switch g1 (w5) @(281,148) /sn:0 /w:[ 0 ] /st:0
  led g5 (.I(w4));   //: @(508,182) /sn:0 /R:3 /w:[ 1 ] /type:0
  FA2 g0 (.A(w5), .B(w6), .Cin(w7), .Cout(w3), .S(w4));   //: @(329, 118) /sz:(137, 126) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 To0<0 Ro0<0 ]

endmodule
