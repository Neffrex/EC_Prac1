//: version "1.8.7"

module CLA16b(B, S, Cout, A, PG, Cin);
//: interface  /sz:(108, 107) /bd:[ Ti0>A[15:0](34/108) Ti1>B[15:0](73/108) Ri0>Cin(53/107) Lo0<Cout(52/107) Bo0<S[15:0](47/108) Bo1<PG(79/108) ]
input [15:0] B;    //: /sn:0 {0}(560,37)(522,37){1}
//: {2}(521,37)(402,37){3}
//: {4}(401,37)(286,37){5}
//: {6}(285,37)(162,37){7}
//: {8}(161,37)(79,37){9}
input [15:0] A;    //: /sn:0 {0}(560,22)(484,22){1}
//: {2}(483,22)(364,22){3}
//: {4}(363,22)(248,22){5}
//: {6}(247,22)(124,22){7}
//: {8}(123,22)(79,22){9}
output PG;    //: /sn:0 {0}(486,302)(486,334){1}
input Cin;    //: /sn:0 {0}(598,92)(598,106){1}
//: {2}(596,108)(550,108){3}
//: {4}(598,110)(598,266)(562,266){5}
output Cout;    //: /sn:0 {0}(74,331)(74,270)(95,270){1}
output [15:0] S;    //: /sn:0 /dp:1 {0}(78,193)(41,193){1}
wire w16;    //: /sn:0 {0}(418,152)(418,235){1}
wire [3:0] w13;    //: /sn:0 {0}(364,63)(364,26){1}
wire [3:0] w6;    //: /sn:0 {0}(286,64)(286,41){1}
wire [3:0] w7;    //: /sn:0 {0}(248,64)(248,26){1}
wire [3:0] w25;    //: /sn:0 /dp:1 {0}(84,188)(266,188)(266,153){1}
wire [3:0] w4;    //: /sn:0 {0}(142,155)(142,178)(84,178){1}
wire w22;    //: /sn:0 /dp:1 {0}(538,151)(538,235){1}
wire w3;    //: /sn:0 {0}(162,155)(162,235){1}
wire [3:0] w0;    //: /sn:0 {0}(162,66)(162,41){1}
wire [3:0] w19;    //: /sn:0 {0}(484,62)(484,26){1}
wire [3:0] w18;    //: /sn:0 {0}(522,62)(522,41){1}
wire [3:0] w12;    //: /sn:0 {0}(402,63)(402,41){1}
wire w23;    //: /sn:0 /dp:1 {0}(522,151)(522,235){1}
wire w10;    //: /sn:0 {0}(302,153)(302,235){1}
wire [3:0] w1;    //: /sn:0 {0}(124,66)(124,26){1}
wire w8;    //: /sn:0 {0}(314,110)(325,110)(325,235){1}
wire w17;    //: /sn:0 {0}(402,152)(402,235){1}
wire w35;    //: /sn:0 {0}(449,235)(449,109)(430,109){1}
wire w33;    //: /sn:0 {0}(201,235)(201,112)(190,112){1}
wire [3:0] w2;    //: /sn:0 /dp:1 {0}(84,208)(502,208)(502,151){1}
wire w11;    //: /sn:0 {0}(286,153)(286,235){1}
wire [3:0] w15;    //: /sn:0 {0}(382,152)(382,198)(84,198){1}
wire w5;    //: /sn:0 {0}(178,155)(178,235){1}
//: enddecls

  //: input g8 (B) @(77,37) /sn:0 /w:[ 9 ]
  Carrylookahead_logic g4 (.P3(w3), .G0(w22), .G1(w16), .G2(w10), .G3(w5), .P0(w23), .P1(w17), .P2(w11), .Cin(Cin), .C1(w35), .C2(w8), .C3(w33), .C4(Cout), .PG(PG));   //: @(96, 236) /sz:(465, 65) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Ri0>5 To0<0 To1<1 To2<0 Lo0<1 Bo0<0 ]
  tran g16(.Z(w0), .I(B[15:12]));   //: @(162,35) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  CLA g3 (.A(w19), .B(w18), .Cin(Cin), .PG(w23), .GG(w22), .S(w2));   //: @(462, 63) /sz:(87, 87) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>3 Bo0<0 Bo1<0 Bo2<1 ]
  //: output g17 (S) @(44,193) /sn:0 /R:2 /w:[ 1 ]
  CLA g2 (.A(w13), .B(w12), .Cin(w35), .PG(w17), .GG(w16), .S(w15));   //: @(342, 64) /sz:(87, 87) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<0 Bo2<0 ]
  CLA g1 (.A(w7), .B(w6), .Cin(w8), .PG(w11), .GG(w10), .S(w25));   //: @(226, 65) /sz:(87, 87) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Bo0<0 Bo1<0 Bo2<1 ]
  concat g18 (.I0(w2), .I1(w15), .I2(w25), .I3(w4), .Z(S));   //: @(79,193) /sn:0 /R:2 /w:[ 0 1 0 1 0 ] /dr:1
  tran g10(.Z(w7), .I(A[11:8]));   //: @(248,20) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  //: output g6 (Cout) @(74,328) /sn:0 /R:3 /w:[ 0 ]
  tran g9(.Z(w1), .I(A[15:12]));   //: @(124,20) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  //: input g7 (A) @(77,22) /sn:0 /w:[ 9 ]
  tran g12(.Z(w19), .I(A[3:0]));   //: @(484,20) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g14(.Z(w12), .I(B[7:4]));   //: @(402,35) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g11(.Z(w13), .I(A[7:4]));   //: @(364,20) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  //: output g5 (PG) @(486,331) /sn:0 /R:3 /w:[ 1 ]
  //: input g19 (Cin) @(598,90) /sn:0 /R:3 /w:[ 0 ]
  //: joint g20 (Cin) @(598, 108) /w:[ -1 1 2 4 ]
  tran g15(.Z(w6), .I(B[11:8]));   //: @(286,35) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  CLA g0 (.A(w1), .B(w0), .Cin(w33), .PG(w3), .GG(w5), .S(w4));   //: @(102, 67) /sz:(87, 87) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<0 Bo2<0 ]
  tran g13(.Z(w18), .I(B[3:0]));   //: @(522,35) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1

endmodule

module PFA(P, S, Cin, B, G, A);
//: interface  /sz:(50, 50) /bd:[ Ti0>A(13/50) Ti1>B(37/50) Ri0>Cin(22/50) Bo0<S(40/50) Bo1<G(25/50) Bo2<P(12/50) ]
input B;    //: /sn:0 {0}(124,181)(135,181){1}
//: {2}(139,181)(184,181){3}
//: {4}(137,183)(137,216){5}
//: {6}(139,218)(212,218){7}
//: {8}(137,220)(137,242)(211,242){9}
input A;    //: /sn:0 {0}(124,171)(143,171){1}
//: {2}(147,171)(174,171)(174,176)(184,176){3}
//: {4}(145,173)(145,211){5}
//: {6}(147,213)(212,213){7}
//: {8}(145,215)(145,237)(211,237){9}
output G;    //: /sn:0 /dp:1 {0}(232,240)(289,240){1}
input Cin;    //: /sn:0 {0}(124,192)(234,192)(234,189)(244,189){1}
output P;    //: /sn:0 /dp:1 {0}(233,216)(288,216){1}
output S;    //: /sn:0 /dp:1 {0}(265,187)(288,187){1}
wire w2;    //: /sn:0 {0}(205,179)(234,179)(234,184)(244,184){1}
//: enddecls

  and g8 (.I0(A), .I1(B), .Z(G));   //: @(222,240) /sn:0 /delay:" 3" /w:[ 9 9 0 ]
  //: output g4 (P) @(285,216) /sn:0 /w:[ 1 ]
  //: output g3 (S) @(285,187) /sn:0 /w:[ 1 ]
  //: input g2 (Cin) @(122,192) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(122,181) /sn:0 /w:[ 0 ]
  //: joint g10 (B) @(137, 181) /w:[ 2 -1 1 4 ]
  xor g6 (.I0(A), .I1(B), .Z(w2));   //: @(195,179) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  or g9 (.I0(A), .I1(B), .Z(P));   //: @(223,216) /sn:0 /delay:" 3" /w:[ 7 7 0 ]
  xor g7 (.I0(w2), .I1(Cin), .Z(S));   //: @(255,187) /sn:0 /delay:" 4" /w:[ 1 1 0 ]
  //: joint g12 (A) @(145, 213) /w:[ 6 5 -1 8 ]
  //: joint g11 (A) @(145, 171) /w:[ 2 -1 1 4 ]
  //: output g5 (G) @(286,240) /sn:0 /w:[ 1 ]
  //: input g0 (A) @(122,171) /sn:0 /w:[ 0 ]
  //: joint g13 (B) @(137, 218) /w:[ 6 5 -1 8 ]

endmodule

module Carrylookahead_logic(P1, C3, G2, P2, G3, C1, P0, G0, C2, G1, Cin, PG, P3, C4);
//: interface  /sz:(312, 40) /bd:[ Ti0>P2(95/312) Ti1>P1(186/312) Ti2>P0(273/312) Ti3>G3(30/312) Ti4>G2(109/312) Ti5>G1(199/312) Ti6>G0(286/312) Ti7>P3(17/312) Ri0>Cin(21/40) To0<C3(71/312) To1<C2(147/312) To2<C1(237/312) Lo0<C4(19/40) Bo0<PG(262/312) ]
input G2;    //: /sn:0 {0}(560,112)(560,172){1}
input P1;    //: /sn:0 {0}(506,114)(506,173){1}
output C3;    //: /sn:0 /dp:1 {0}(287,338)(287,374){1}
output PG;    //: /sn:0 /dp:1 {0}(26,258)(26,261){1}
//: {2}(28,263)(47,263)(47,272){3}
//: {4}(26,265)(26,383){5}
input G0;    //: /sn:0 {0}(580,112)(580,172){1}
output C4;    //: /sn:0 /dp:1 {0}(112,383)(112,336){1}
output C2;    //: /sn:0 /dp:1 {0}(403,336)(403,373){1}
input Cin;    //: /sn:0 {0}(582,233)(471,233){1}
//: {2}(467,233)(381,233){3}
//: {4}(377,233)(239,233){5}
//: {6}(235,233)(52,233)(52,272){7}
//: {8}(237,235)(237,257){9}
//: {10}(379,235)(379,262){11}
//: {12}(469,235)(469,248){13}
input P3;    //: /sn:0 {0}(486,113)(486,173){1}
input G1;    //: /sn:0 {0}(570,112)(570,172){1}
input G3;    //: /sn:0 {0}(550,112)(550,172){1}
input P0;    //: /sn:0 {0}(516,113)(516,173){1}
output C1;    //: /sn:0 {0}(484,373)(484,338){1}
input P2;    //: /sn:0 {0}(496,114)(496,173){1}
wire w6;    //: /sn:0 {0}(374,283)(374,305)(398,305)(398,315){1}
wire [3:0] w13;    //: /sn:0 {0}(-6,205)(17,205){1}
//: {2}(18,205)(22,205){3}
//: {4}(23,205)(27,205){5}
//: {6}(28,205)(32,205){7}
//: {8}(33,205)(78,205){9}
//: {10}(79,205)(83,205){11}
//: {12}(84,205)(88,205){13}
//: {14}(89,205)(117,205){15}
//: {16}(118,205)(122,205){17}
//: {18}(123,205)(157,205){19}
//: {20}(158,205)(264,205){21}
//: {22}(265,205)(269,205){23}
//: {24}(270,205)(307,205){25}
//: {26}(308,205)(368,205){27}
//: {28}(369,205)(373,205){29}
//: {30}(374,205)(399,205){31}
//: {32}(400,205)(463,205){33}
//: {34}(464,205)(501,205)(501,179){35}
wire [3:0] w16;    //: /sn:0 {0}(20,216)(93,216){1}
//: {2}(94,216)(127,216){3}
//: {4}(128,216)(162,216){5}
//: {6}(163,216)(186,216){7}
//: {8}(187,216)(221,216){9}
//: {10}(222,216)(226,216){11}
//: {12}(227,216)(231,216){13}
//: {14}(232,216)(274,216){15}
//: {16}(275,216)(312,216){17}
//: {18}(313,216)(338,216){19}
//: {20}(339,216)(404,216){21}
//: {22}(405,216)(434,216){23}
//: {24}(435,216)(485,216){25}
//: {26}(486,216)(565,216)(565,178){27}
wire w7;    //: /sn:0 {0}(313,220)(313,258){1}
wire w34;    //: /sn:0 {0}(123,276)(123,297)(112,297)(112,315){1}
wire w4;    //: /sn:0 {0}(308,209)(308,258){1}
wire w25;    //: /sn:0 {0}(128,220)(128,255){1}
wire w0;    //: /sn:0 {0}(400,209)(400,264){1}
wire w22;    //: /sn:0 {0}(464,209)(464,248){1}
wire w3;    //: /sn:0 {0}(486,220)(486,317){1}
wire w36;    //: /sn:0 {0}(89,209)(89,255){1}
wire w30;    //: /sn:0 {0}(232,220)(232,257){1}
wire w29;    //: /sn:0 {0}(123,209)(123,255){1}
wire w37;    //: /sn:0 {0}(87,276)(87,302)(107,302)(107,315){1}
wire w42;    //: /sn:0 {0}(84,255)(84,209){1}
wire w19;    //: /sn:0 {0}(28,209)(28,237){1}
wire w18;    //: /sn:0 {0}(33,209)(33,237){1}
wire w12;    //: /sn:0 {0}(405,220)(405,264){1}
wire w23;    //: /sn:0 {0}(23,237)(23,209){1}
wire w10;    //: /sn:0 {0}(275,220)(275,256){1}
wire w21;    //: /sn:0 {0}(435,220)(435,300)(408,300)(408,315){1}
wire w24;    //: /sn:0 {0}(161,277)(161,302)(117,302)(117,315){1}
wire w1;    //: /sn:0 {0}(369,262)(369,209){1}
wire w31;    //: /sn:0 {0}(230,278)(230,308)(279,308)(279,317){1}
wire w32;    //: /sn:0 {0}(227,257)(227,220){1}
wire w8;    //: /sn:0 {0}(311,279)(311,303)(289,303)(289,317){1}
wire w17;    //: /sn:0 {0}(187,220)(187,305)(122,305)(122,315){1}
wire w27;    //: /sn:0 {0}(467,269)(467,300)(481,300)(481,317){1}
wire w28;    //: /sn:0 {0}(270,277)(270,303)(284,303)(284,317){1}
wire w33;    //: /sn:0 {0}(222,257)(222,220){1}
wire w35;    //: /sn:0 {0}(94,220)(94,255){1}
wire w45;    //: /sn:0 {0}(50,293)(50,310)(102,310)(102,315){1}
wire w14;    //: /sn:0 {0}(158,209)(158,256){1}
wire w11;    //: /sn:0 {0}(339,220)(339,308)(294,308)(294,317){1}
wire w2;    //: /sn:0 {0}(265,256)(265,209){1}
wire w41;    //: /sn:0 {0}(118,255)(118,209){1}
wire w15;    //: /sn:0 {0}(163,220)(163,256){1}
wire w38;    //: /sn:0 {0}(18,237)(18,209){1}
wire w5;    //: /sn:0 {0}(374,209)(374,262){1}
wire w43;    //: /sn:0 {0}(79,255)(79,209){1}
wire w9;    //: /sn:0 {0}(403,285)(403,315){1}
wire w26;    //: /sn:0 {0}(270,209)(270,256){1}
//: enddecls

  //: input g4 (P1) @(506,112) /sn:0 /R:3 /w:[ 0 ]
  //: output g8 (C3) @(287,371) /sn:0 /R:3 /w:[ 1 ]
  //: joint g44 (Cin) @(237, 233) /w:[ 5 -1 6 8 ]
  //: input g3 (G2) @(560,110) /sn:0 /R:3 /w:[ 0 ]
  and g16 (.I0(Cin), .I1(w5), .I2(w1), .Z(w6));   //: @(374,273) /sn:0 /R:3 /delay:" 3" /w:[ 11 1 0 0 ]
  and g47 (.I0(w35), .I1(w36), .I2(w42), .I3(w43), .Z(w37));   //: @(87,266) /sn:0 /R:3 /delay:" 3" /w:[ 1 1 0 0 0 ]
  and g17 (.I0(w0), .I1(w12), .Z(w9));   //: @(403,275) /sn:0 /R:3 /delay:" 3" /w:[ 1 1 0 ]
  tran g26(.Z(w11), .I(w16[2]));   //: @(339,214) /sn:0 /R:1 /w:[ 0 19 20 ] /ss:1
  //: input g2 (P2) @(496,112) /sn:0 /R:3 /w:[ 0 ]
  tran g23(.Z(w21), .I(w16[1]));   //: @(435,214) /sn:0 /R:1 /w:[ 0 23 24 ] /ss:1
  tran g30(.Z(w1), .I(w13[1]));   //: @(369,203) /sn:0 /R:1 /w:[ 1 27 28 ] /ss:1
  //: input g1 (G3) @(550,110) /sn:0 /R:3 /w:[ 0 ]
  or g24 (.I0(w11), .I1(w8), .I2(w28), .I3(w31), .Z(C3));   //: @(287,328) /sn:0 /R:3 /delay:" 3" /w:[ 1 1 1 1 0 ]
  tran g39(.Z(w26), .I(w13[1]));   //: @(270,203) /sn:0 /R:1 /w:[ 0 23 24 ] /ss:1
  tran g29(.Z(w12), .I(w16[0]));   //: @(405,214) /sn:0 /R:1 /w:[ 0 21 22 ] /ss:1
  tran g51(.Z(w25), .I(w16[1]));   //: @(128,214) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  tran g18(.Z(w22), .I(w13[0]));   //: @(464,203) /sn:0 /R:1 /w:[ 0 33 34 ] /ss:1
  tran g65(.Z(w38), .I(w13[3]));   //: @(18,203) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: output g10 (C1) @(484,370) /sn:0 /R:3 /w:[ 0 ]
  or g25 (.I0(w17), .I1(w24), .I2(w34), .I3(w37), .I4(w45), .Z(C4));   //: @(112,326) /sn:0 /R:3 /delay:" 3" /w:[ 1 1 1 1 1 1 ]
  and g64 (.I0(w18), .I1(w19), .I2(w23), .I3(w38), .Z(PG));   //: @(26,248) /sn:0 /R:3 /delay:" 3" /w:[ 1 1 0 0 0 ]
  tran g49(.Z(w14), .I(w13[3]));   //: @(158,203) /sn:0 /R:1 /w:[ 0 19 20 ] /ss:1
  //: input g6 (P0) @(516,111) /sn:0 /R:3 /w:[ 0 ]
  tran g50(.Z(w15), .I(w16[2]));   //: @(163,214) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: joint g58 (PG) @(26, 263) /w:[ 2 1 -1 4 ]
  tran g68(.Z(w18), .I(w13[0]));   //: @(33,203) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  //: input g7 (G0) @(580,110) /sn:0 /R:3 /w:[ 0 ]
  //: output g9 (C2) @(403,370) /sn:0 /R:3 /w:[ 1 ]
  and g35 (.I0(Cin), .I1(w30), .I2(w32), .I3(w33), .Z(w31));   //: @(230,268) /sn:0 /R:3 /delay:" 3" /w:[ 9 1 0 0 0 ]
  tran g56(.Z(w42), .I(w13[2]));   //: @(84,203) /sn:0 /R:1 /w:[ 1 11 12 ] /ss:1
  concat g22 (.I0(G0), .I1(G1), .I2(G2), .I3(G3), .Z(w16));   //: @(565,177) /sn:0 /R:3 /w:[ 1 1 1 1 27 ] /dr:1
  tran g31(.Z(w5), .I(w13[0]));   //: @(374,203) /sn:0 /R:1 /w:[ 0 29 30 ] /ss:1
  tran g67(.Z(w19), .I(w13[1]));   //: @(28,203) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  and g33 (.I0(w4), .I1(w7), .Z(w8));   //: @(311,269) /sn:0 /R:3 /delay:" 3" /w:[ 1 1 0 ]
  tran g36(.Z(w4), .I(w13[2]));   //: @(308,203) /sn:0 /R:1 /w:[ 0 25 26 ] /ss:1
  tran g41(.Z(w33), .I(w16[2]));   //: @(222,214) /sn:0 /R:1 /w:[ 1 9 10 ] /ss:1
  and g45 (.I0(w14), .I1(w15), .Z(w24));   //: @(161,267) /sn:0 /R:3 /delay:" 3" /w:[ 1 1 0 ]
  tran g54(.Z(w35), .I(w16[0]));   //: @(94,214) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g40(.Z(w10), .I(w16[0]));   //: @(275,214) /sn:0 /R:1 /w:[ 0 15 16 ] /ss:1
  tran g42(.Z(w32), .I(w16[1]));   //: @(227,214) /sn:0 /R:1 /w:[ 1 11 12 ] /ss:1
  tran g52(.Z(w29), .I(w13[2]));   //: @(123,203) /sn:0 /R:1 /w:[ 0 17 18 ] /ss:1
  tran g66(.Z(w23), .I(w13[2]));   //: @(23,203) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  and g12 (.I0(w22), .I1(Cin), .Z(w27));   //: @(467,259) /sn:0 /R:3 /delay:" 3" /w:[ 1 13 0 ]
  tran g28(.Z(w0), .I(w13[1]));   //: @(400,203) /sn:0 /R:1 /w:[ 0 31 32 ] /ss:1
  and g34 (.I0(w10), .I1(w26), .I2(w2), .Z(w28));   //: @(270,267) /sn:0 /R:3 /delay:" 3" /w:[ 1 1 0 0 ]
  and g46 (.I0(w25), .I1(w29), .I2(w41), .Z(w34));   //: @(123,266) /sn:0 /R:3 /delay:" 3" /w:[ 1 1 0 0 ]
  tran g57(.Z(w43), .I(w13[3]));   //: @(79,203) /sn:0 /R:1 /w:[ 1 9 10 ] /ss:1
  //: input g5 (G1) @(570,110) /sn:0 /R:3 /w:[ 0 ]
  or g11 (.I0(w27), .I1(w3), .Z(C1));   //: @(484,328) /sn:0 /R:3 /delay:" 3" /w:[ 1 1 1 ]
  //: input g14 (Cin) @(584,233) /sn:0 /R:2 /w:[ 0 ]
  concat g21 (.I0(P0), .I1(P1), .I2(P2), .I3(P3), .Z(w13));   //: @(501,178) /sn:0 /R:3 /w:[ 1 1 1 1 35 ] /dr:1
  //: joint g19 (Cin) @(469, 233) /w:[ 1 -1 2 12 ]
  tran g20(.Z(w3), .I(w16[0]));   //: @(486,214) /sn:0 /R:1 /w:[ 0 25 26 ] /ss:1
  //: joint g32 (Cin) @(379, 233) /w:[ 3 -1 4 10 ]
  //: output g63 (PG) @(26,380) /sn:0 /R:3 /w:[ 5 ]
  //: input g0 (P3) @(486,111) /sn:0 /R:3 /w:[ 0 ]
  or g15 (.I0(w21), .I1(w9), .I2(w6), .Z(C2));   //: @(403,326) /sn:0 /R:3 /delay:" 3" /w:[ 1 1 1 0 ]
  tran g38(.Z(w2), .I(w13[2]));   //: @(265,203) /sn:0 /R:1 /w:[ 1 21 22 ] /ss:1
  tran g43(.Z(w30), .I(w16[0]));   //: @(232,214) /sn:0 /R:1 /w:[ 0 13 14 ] /ss:1
  and g48 (.I0(PG), .I1(Cin), .Z(w45));   //: @(50,283) /sn:0 /R:3 /delay:" 3" /w:[ 3 7 0 ]
  tran g27(.Z(w17), .I(w16[3]));   //: @(187,214) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g37(.Z(w7), .I(w16[1]));   //: @(313,214) /sn:0 /R:1 /w:[ 0 17 18 ] /ss:1
  tran g55(.Z(w36), .I(w13[1]));   //: @(89,203) /sn:0 /R:1 /w:[ 0 13 14 ] /ss:1
  //: output g13 (C4) @(112,380) /sn:0 /R:3 /w:[ 0 ]
  tran g53(.Z(w41), .I(w13[3]));   //: @(118,203) /sn:0 /R:1 /w:[ 1 15 16 ] /ss:1

endmodule

module main;    //: root_module
wire [15:0] w6;    //: /sn:0 /dp:1 {0}(226,96)(226,129)(289,129)(289,139){1}
wire [15:0] w7;    //: /sn:0 {0}(394,93)(394,127)(328,127)(328,139){1}
wire w0;    //: /sn:0 {0}(395,193)(364,193){1}
wire w2;    //: /sn:0 {0}(254,192)(218,192){1}
wire w5;    //: /sn:0 {0}(334,248)(334,278)(356,278){1}
wire [15:0] w9;    //: /sn:0 {0}(322,361)(302,361)(302,360){1}
//: {2}(302,356)(302,317){3}
//: {4}(304,315)(350,315){5}
//: {6}(302,313)(302,248){7}
//: {8}(300,358)(253,358){9}
//: enddecls

  //: switch g8 (w0) @(413,193) /sn:0 /R:2 /w:[ 0 ] /st:0
  led g4 (.I(w5));   //: @(363,278) /sn:0 /R:3 /w:[ 1 ] /type:0
  led g3 (.I(w2));   //: @(211,192) /sn:0 /R:1 /w:[ 1 ] /type:0
  //: dip g2 (w7) @(394,83) /sn:0 /w:[ 0 ] /st:16
  //: dip g1 (w6) @(226,86) /sn:0 /w:[ 0 ] /st:16
  //: joint g10 (w9) @(302, 358) /w:[ -1 2 8 1 ]
  led g6 (.I(w9));   //: @(329,361) /sn:0 /R:3 /w:[ 0 ] /type:3
  led g9 (.I(w9));   //: @(246,358) /sn:0 /R:1 /w:[ 9 ] /type:2
  //: joint g7 (w9) @(302, 315) /w:[ 4 6 -1 3 ]
  led g5 (.I(w9));   //: @(357,315) /sn:0 /R:3 /w:[ 5 ] /type:1
  CLA16b g0 (.B(w7), .A(w6), .Cin(w0), .Cout(w2), .PG(w5), .S(w9));   //: @(255, 140) /sz:(108, 107) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 Bo1<7 ]

endmodule

module CLA(A, S, GG, Cin, PG, B);
//: interface  /sz:(87, 87) /bd:[ Ti0>B[3:0](60/87) Ti1>A[3:0](22/87) Ri0>Cin(45/87) Bo0<S[3:0](40/87) Bo1<GG(76/87) Bo2<PG(60/87) ]
input [3:0] B;    //: /sn:0 {0}(140,107)(193,107){1}
//: {2}(194,107)(285,107){3}
//: {4}(286,107)(383,107){5}
//: {6}(384,107)(477,107){7}
//: {8}(478,107)(492,107){9}
output GG;    //: /sn:0 {0}(151,283)(114,283)(114,321){1}
input [3:0] A;    //: /sn:0 {0}(141,91)(169,91){1}
//: {2}(170,91)(261,91){3}
//: {4}(262,91)(359,91){5}
//: {6}(360,91)(453,91){7}
//: {8}(454,91)(490,91){9}
output PG;    //: /sn:0 {0}(414,336)(414,302){1}
input Cin;    //: /sn:0 /dp:1 {0}(464,167)(504,167){1}
//: {2}(506,165)(506,101)(528,101){3}
//: {4}(506,169)(506,282)(465,282){5}
output [3:0] S;    //: /sn:0 {0}(84,230)(129,230){1}
wire w6;    //: /sn:0 {0}(274,145)(274,127)(286,127)(286,111){1}
wire w13;    //: /sn:0 {0}(339,145)(339,119)(360,119)(360,95){1}
wire w16;    //: /sn:0 {0}(351,197)(351,260){1}
wire w7;    //: /sn:0 {0}(248,145)(248,119)(262,119)(262,95){1}
wire w4;    //: /sn:0 {0}(182,194)(182,260){1}
wire w39;    //: /sn:0 /dp:1 {0}(389,260)(389,168)(377,168){1}
wire w0;    //: /sn:0 {0}(194,142)(194,111){1}
wire w37;    //: /sn:0 /dp:1 {0}(223,260)(223,165)(208,165){1}
wire w12;    //: /sn:0 {0}(363,145)(363,127)(384,127)(384,111){1}
wire w18;    //: /sn:0 {0}(450,144)(450,124)(478,124)(478,111){1}
wire w19;    //: /sn:0 {0}(426,144)(426,116)(454,116)(454,95){1}
wire w10;    //: /sn:0 {0}(261,200)(261,260){1}
wire w23;    //: /sn:0 {0}(453,196)(453,215)(135,215){1}
wire w24;    //: /sn:0 /dp:1 {0}(277,200)(277,235)(135,235){1}
wire w1;    //: /sn:0 {0}(170,142)(170,95){1}
wire w46;    //: /sn:0 {0}(338,197)(338,260){1}
wire w17;    //: /sn:0 {0}(366,197)(366,225)(135,225){1}
wire w27;    //: /sn:0 /dp:1 {0}(425,260)(425,196){1}
wire w33;    //: /sn:0 /dp:1 {0}(438,260)(438,196){1}
wire w5;    //: /sn:0 {0}(197,194)(197,245)(135,245){1}
wire w38;    //: /sn:0 /dp:1 {0}(299,260)(299,170)(289,170){1}
wire w9;    //: /sn:0 {0}(247,200)(247,260){1}
wire w26;    //: /sn:0 {0}(169,194)(169,260){1}
//: enddecls

  //: input g4 (A) @(139,91) /sn:0 /w:[ 0 ]
  //: output g8 (S) @(87,230) /sn:0 /R:2 /w:[ 0 ]
  PFA g3 (.A(w19), .B(w18), .Cin(Cin), .S(w23), .G(w33), .P(w27));   //: @(413, 145) /sz:(50, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Bo0<0 Bo1<1 Bo2<1 ]
  tran g16(.Z(w0), .I(B[3]));   //: @(194,105) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: joint g17 (Cin) @(506, 167) /w:[ -1 2 1 4 ]
  PFA g2 (.A(w13), .B(w12), .Cin(w39), .S(w17), .G(w16), .P(w46));   //: @(326, 146) /sz:(50, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<0 Bo2<0 ]
  Carrylookahead_logic g30 (.P3(w26), .G0(w33), .G1(w16), .G2(w10), .G3(w4), .P0(w27), .P1(w46), .P2(w9), .Cin(Cin), .C1(w39), .C2(w38), .C3(w37), .C4(GG), .PG(PG));   //: @(152, 261) /sz:(312, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>1 Ti3>1 Ti4>1 Ti5>0 Ti6>1 Ti7>1 Ri0>5 To0<0 To1<0 To2<0 Lo0<0 Bo0<1 ]
  PFA g1 (.A(w7), .B(w6), .Cin(w38), .S(w24), .G(w10), .P(w9));   //: @(234, 146) /sz:(54, 53) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<0 Bo2<0 ]
  concat g29 (.I0(w23), .I1(w17), .I2(w24), .I3(w5), .Z(S));   //: @(130,230) /sn:0 /R:2 /w:[ 1 1 1 1 1 ] /dr:0
  //: output g18 (GG) @(114,318) /sn:0 /R:3 /w:[ 1 ]
  tran g10(.Z(w13), .I(A[1]));   //: @(360,89) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g6 (Cin) @(530,101) /sn:0 /R:2 /w:[ 3 ]
  //: output g7 (PG) @(414,333) /sn:0 /R:3 /w:[ 0 ]
  tran g9(.Z(w19), .I(A[0]));   //: @(454,89) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g12(.Z(w1), .I(A[3]));   //: @(170,89) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: input g5 (B) @(138,107) /sn:0 /w:[ 0 ]
  tran g11(.Z(w7), .I(A[2]));   //: @(262,89) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g14(.Z(w12), .I(B[1]));   //: @(384,105) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  PFA g0 (.A(w1), .B(w0), .Cin(w37), .S(w5), .G(w4), .P(w26));   //: @(157, 143) /sz:(50, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<0 Bo2<0 ]
  tran g15(.Z(w6), .I(B[2]));   //: @(286,105) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g13(.Z(w18), .I(B[0]));   //: @(478,105) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1

endmodule
