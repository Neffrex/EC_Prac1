//: version "1.8.7"

module HA(C, S, B, A);
//: interface  /sz:(263, 230) /bd:[ Li0>A(49/230) Li1>B(127/230) To0<C(143/263) Ro0<S(91/230) ]
input B;    //: /sn:0 {0}(122,340)(208,340){1}
//: {2}(212,340)(257,340)(257,326)(265,326){3}
//: {4}(210,342)(210,371)(265,371){5}
input A;    //: /sn:0 {0}(122,321)(225,321){1}
//: {2}(229,321)(265,321){3}
//: {4}(227,323)(227,366)(265,366){5}
output C;    //: /sn:0 /dp:1 {0}(286,369)(380,369){1}
output S;    //: /sn:0 /dp:1 {0}(286,324)(375,324){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(276,324) /sn:0 /delay:" 5" /w:[ 3 3 0 ]
  //: output g3 (C) @(377,369) /sn:0 /w:[ 1 ]
  //: output g2 (S) @(372,324) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(120,340) /sn:0 /w:[ 0 ]
  //: joint g6 (B) @(210, 340) /w:[ 2 -1 1 4 ]
  //: joint g7 (A) @(227, 321) /w:[ 2 -1 1 4 ]
  and g5 (.I0(A), .I1(B), .Z(C));   //: @(276,369) /sn:0 /delay:" 4" /w:[ 5 5 0 ]
  //: input g0 (A) @(120,321) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(206,191)(265,191){1}
wire w7;    //: /sn:0 {0}(208,233)(265,233){1}
wire w4;    //: /sn:0 {0}(436,190)(472,190){1}
wire w3;    //: /sn:0 {0}(364,106)(364,76){1}
wire w5;    //: /sn:0 {0}(206,150)(265,150){1}
//: enddecls

  led g4 (.I(w3));   //: @(364,69) /sn:0 /w:[ 1 ] /type:0
  //: switch g3 (w7) @(191,233) /sn:0 /w:[ 0 ] /st:0
  //: switch g2 (w6) @(189,191) /sn:0 /w:[ 0 ] /st:1
  //: switch g1 (w5) @(189,150) /sn:0 /w:[ 0 ] /st:0
  led g5 (.I(w4));   //: @(479,190) /sn:0 /R:3 /w:[ 1 ] /type:0
  FA g0 (.A(w5), .B(w6), .Cin(w7), .Cout(w3), .S(w4));   //: @(266, 107) /sz:(169, 168) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 To0<0 Ro0<0 ]

endmodule

module FA(Cout, S, Cin, B, A);
//: interface  /sz:(169, 168) /bd:[ Li0>A(43/168) Li1>B(84/168) Li2>Cin(126/168) To0<Cout(98/169) Ro0<S(83/168) ]
input B;    //: /sn:0 {0}(125,198)(216,198){1}
input A;    //: /sn:0 {0}(125,181)(216,181){1}
input Cin;    //: /sn:0 {0}(132,107)(277,107){1}
output Cout;    //: /sn:0 /dp:1 {0}(391,153)(419,153){1}
output S;    //: /sn:0 {0}(299,98)(299,67)(317,67){1}
wire w1;    //: /sn:0 {0}(239,175)(239,155)(370,155){1}
wire w8;    //: /sn:0 {0}(259,199)(269,199)(269,121)(277,121){1}
wire w5;    //: /sn:0 {0}(319,114)(360,114)(360,150)(370,150){1}
//: enddecls

  //: output g4 (Cout) @(416,153) /sn:0 /w:[ 1 ]
  //: output g3 (S) @(314,67) /sn:0 /w:[ 1 ]
  //: input g2 (Cin) @(130,107) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(123,198) /sn:0 /w:[ 0 ]
  HA g6 (.B(w8), .A(Cin), .S(S), .C(w5));   //: @(278, 99) /sz:(40, 40) /sn:0 /p:[ Li0>1 Li1>1 To0<0 Ro0<0 ]
  or g9 (.I0(w5), .I1(w1), .Z(Cout));   //: @(381,153) /sn:0 /delay:" 4" /w:[ 1 1 0 ]
  HA g5 (.B(B), .A(A), .C(w1), .S(w8));   //: @(217, 176) /sz:(41, 40) /sn:0 /p:[ Li0>1 Li1>1 To0<0 Ro0<0 ]
  //: input g0 (A) @(123,181) /sn:0 /w:[ 0 ]

endmodule
