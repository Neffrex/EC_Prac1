//: version "1.8.7"

module FA2(Cout, S, Cin, B, A);
//: interface  /sz:(137, 126) /bd:[ Li0>A(30/126) Li1>B(66/126) Li2>Cin(101/126) To0<Cout(72/137) Ro0<S(64/126) ]
input B;    //: /sn:0 {0}(144,181)(144,255){1}
//: {2}(146,257)(218,257){3}
//: {4}(144,259)(144,377){5}
//: {6}(146,379)(159,379)(159,376)(218,376){7}
//: {8}(144,381)(144,415)(218,415){9}
input A;    //: /sn:0 {0}(113,181)(113,239){1}
//: {2}(115,241)(208,241)(208,252)(218,252){3}
//: {4}(113,243)(113,312){5}
//: {6}(115,314)(126,314)(126,323)(219,323){7}
//: {8}(113,316)(113,371)(218,371){9}
input Cin;    //: /sn:0 {0}(173,180)(173,270){1}
//: {2}(175,272)(341,272){3}
//: {4}(173,274)(173,326){5}
//: {6}(175,328)(219,328){7}
//: {8}(173,330)(173,420)(218,420){9}
output Cout;    //: /sn:0 {0}(392,381)(455,381){1}
output S;    //: /sn:0 {0}(362,270)(451,270){1}
wire w8;    //: /sn:0 {0}(240,326)(280,326)(280,337)(325,337){1}
wire w17;    //: /sn:0 {0}(346,340)(361,340)(361,378)(371,378){1}
wire w14;    //: /sn:0 {0}(239,418)(361,418)(361,383)(371,383){1}
wire w11;    //: /sn:0 {0}(239,374)(283,374)(283,342)(325,342){1}
wire w2;    //: /sn:0 {0}(239,255)(331,255)(331,267)(341,267){1}
//: enddecls

  or g8 (.I0(w8), .I1(w11), .Z(w17));   //: @(336,340) /sn:0 /delay:" 4" /w:[ 1 1 0 ]
  xor g4 (.I0(w2), .I1(Cin), .Z(S));   //: @(352,270) /sn:0 /delay:" 5" /w:[ 1 3 0 ]
  //: output g16 (Cout) @(452,381) /sn:0 /w:[ 1 ]
  xor g3 (.I0(A), .I1(B), .Z(w2));   //: @(229,255) /sn:0 /delay:" 5" /w:[ 3 3 0 ]
  //: output g17 (S) @(448,270) /sn:0 /w:[ 1 ]
  //: input g2 (Cin) @(173,178) /sn:0 /R:3 /w:[ 0 ]
  //: input g1 (B) @(144,179) /sn:0 /R:3 /w:[ 0 ]
  //: joint g10 (B) @(144, 379) /w:[ 6 5 -1 8 ]
  and g6 (.I0(A), .I1(B), .Z(w11));   //: @(229,374) /sn:0 /delay:" 4" /w:[ 9 7 0 ]
  or g9 (.I0(w17), .I1(w14), .Z(Cout));   //: @(382,381) /sn:0 /delay:" 4" /w:[ 1 1 0 ]
  and g7 (.I0(B), .I1(Cin), .Z(w14));   //: @(229,418) /sn:0 /delay:" 4" /w:[ 9 9 0 ]
  //: joint g12 (A) @(113, 314) /w:[ 6 5 -1 8 ]
  //: joint g14 (B) @(144, 257) /w:[ 2 1 -1 4 ]
  //: joint g11 (Cin) @(173, 328) /w:[ 6 5 -1 8 ]
  and g5 (.I0(A), .I1(Cin), .Z(w8));   //: @(230,326) /sn:0 /delay:" 4" /w:[ 7 7 0 ]
  //: joint g15 (Cin) @(173, 272) /w:[ 2 1 -1 4 ]
  //: input g0 (A) @(113,179) /sn:0 /R:3 /w:[ 0 ]
  //: joint g13 (A) @(113, 241) /w:[ 2 1 -1 4 ]

endmodule

module CPA(Cin, B, S, A, Cout);
//: interface  /sz:(327, 51) /bd:[ Ti0>A(106/327) Ti1>B(174/327) Ri0>Cin(24/51) Lo0<C4(28/51) Bo0<S3(44/327) Bo1<S2(118/327) Bo2<S1(203/327) Bo3<S0(280/327) ]
input [3:0] B;    //: /sn:0 {0}(734,44)(698,44){1}
//: {2}(697,44)(597,44){3}
//: {4}(596,44)(500,44){5}
//: {6}(499,44)(399,44){7}
//: {8}(398,44)(319,44){9}
input [3:0] A;    //: /sn:0 {0}(319,21)(377,21){1}
//: {2}(378,21)(471,21){3}
//: {4}(472,21)(572,21){5}
//: {6}(573,21)(671,21){7}
//: {8}(672,21)(725,21){9}
input Cin;    //: /sn:0 /dp:1 {0}(722,125)(749,125){1}
output Cout;    //: /sn:0 /dp:1 {0}(354,113)(331,113)(331,181){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(256,247)(168,247){1}
wire A0;    //: /sn:0 {0}(675,86)(675,33)(672,33)(672,25){1}
wire w6;    //: /sn:0 {0}(500,48)(500,56)(497,56)(497,80){1}
wire w7;    //: /sn:0 {0}(573,25)(573,83){1}
wire S1;    //: /sn:0 {0}(587,155)(587,242)(262,242){1}
wire w4;    //: /sn:0 {0}(620,122)(652,122){1}
wire A3;    //: /sn:0 {0}(377,77)(377,33)(378,33)(378,25){1}
wire w3;    //: /sn:0 {0}(424,116)(450,116){1}
wire w1;    //: /sn:0 /dp:1 {0}(391,149)(391,262)(262,262){1}
wire w8;    //: /sn:0 {0}(597,48)(597,83){1}
wire w2;    //: /sn:0 {0}(472,25)(472,33)(473,33)(473,80){1}
wire B3;    //: /sn:0 {0}(401,77)(401,56)(399,56)(399,48){1}
wire w5;    //: /sn:0 {0}(550,119)(520,119){1}
wire B0;    //: /sn:0 {0}(699,86)(699,56)(698,56)(698,48){1}
wire w9;    //: /sn:0 {0}(689,158)(689,232)(262,232){1}
wire S2;    //: /sn:0 {0}(487,152)(487,252)(262,252){1}
//: enddecls

  //: input g8 (Cin) @(751,125) /sn:0 /R:2 /w:[ 1 ]
  tran g4(.Z(w2), .I(A[2]));   //: @(472,19) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  FA2 g16 (.B(w6), .A(w2), .Cin(w5), .Cout(w3), .S(S2));   //: @(451, 81) /sz:(68, 70) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<0 ]
  tran g3(.Z(w7), .I(A[1]));   //: @(573,19) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  FA2 g17 (.B(B3), .A(A3), .Cin(w3), .Cout(Cout), .S(w1));   //: @(355, 78) /sz:(68, 70) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<0 Bo0<0 ]
  tran g2(.Z(A0), .I(A[0]));   //: @(672,19) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: input g1 (B) @(317,44) /sn:0 /w:[ 9 ]
  tran g18(.Z(w8), .I(B[1]));   //: @(597,42) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  concat g10 (.I0(w9), .I1(S1), .I2(S2), .I3(w1), .Z(S));   //: @(257,247) /sn:0 /R:2 /w:[ 1 1 1 1 0 ] /dr:0
  tran g6(.Z(B3), .I(B[3]));   //: @(399,42) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  //: output g9 (S) @(171,247) /sn:0 /R:2 /w:[ 1 ]
  tran g7(.Z(w6), .I(B[2]));   //: @(500,42) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  FA2 g14 (.B(B0), .A(A0), .Cin(Cin), .Cout(w4), .S(w9));   //: @(653, 87) /sz:(68, 70) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  tran g5(.Z(A3), .I(A[3]));   //: @(378,19) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g19(.Z(B0), .I(B[0]));   //: @(698,42) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  FA2 g15 (.B(w8), .A(w7), .Cin(w4), .Cout(w5), .S(S1));   //: @(551, 84) /sz:(68, 70) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  //: input g0 (A) @(317,21) /sn:0 /w:[ 0 ]
  //: output g13 (Cout) @(331,178) /sn:0 /R:3 /w:[ 1 ]

endmodule

module main;    //: root_module
wire w7;    //: /sn:0 {0}(-9482,-375)(-9492,-375){1}
wire w3;    //: /sn:0 /dp:1 {0}(439,368)(308,368)(308,207)(325,207){1}
wire [3:0] w0;    //: /sn:0 /dp:1 {0}(609,81)(609,145){1}
wire [3:0] w1;    //: /sn:0 /dp:1 {0}(439,378)(396,378)(396,287)(521,287)(521,272){1}
wire w8;    //: /sn:0 /dp:1 {0}(737,206)(768,206){1}
wire w14;    //: /sn:0 {0}(10636,658)(10636,668){1}
wire [3:0] w2;    //: /sn:0 /dp:1 {0}(437,80)(437,145){1}
wire [4:0] w5;    //: /sn:0 {0}(554,350)(554,373)(445,373){1}
//: enddecls

  //: dip g4 (w0) @(609,71) /sn:0 /w:[ 0 ] /st:10
  //: dip g3 (w2) @(437,70) /sn:0 /w:[ 0 ] /st:10
  //: switch g16 (w8) @(786,206) /sn:0 /R:2 /w:[ 1 ] /st:0
  led g2 (.I(w5));   //: @(554,343) /sn:0 /w:[ 0 ] /type:3
  concat g1 (.I0(w1), .I1(w3), .Z(w5));   //: @(444,373) /sn:0 /w:[ 0 0 1 ] /dr:0
  //: switch g6 (w14) @(10636,645) /sn:0 /R:3 /w:[ 0 ] /st:0
  CPA g0 (.B(w0), .A(w2), .Cin(w8), .Cout(w3), .S(w1));   //: @(326, 146) /sz:(410, 125) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  //: switch g15 (w7) @(-9464,-375) /sn:0 /R:2 /w:[ 0 ] /st:0

endmodule
