//: version "1.8.7"

module HA(C, S, B, A);
//: interface  /sz:(263, 230) /bd:[ Li0>B(127/230) Li1>A(49/230) To0<C(143/263) Ro0<S(91/230) ]
input B;    //: /sn:0 {0}(122,340)(208,340){1}
//: {2}(212,340)(257,340)(257,326)(265,326){3}
//: {4}(210,342)(210,371)(265,371){5}
input A;    //: /sn:0 {0}(122,321)(225,321){1}
//: {2}(229,321)(265,321){3}
//: {4}(227,323)(227,366)(265,366){5}
output C;    //: /sn:0 /dp:1 {0}(286,369)(380,369){1}
output S;    //: /sn:0 /dp:1 {0}(286,324)(375,324){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(276,324) /sn:0 /delay:" 5" /w:[ 3 3 0 ]
  //: output g3 (C) @(377,369) /sn:0 /w:[ 1 ]
  //: output g2 (S) @(372,324) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(120,340) /sn:0 /w:[ 0 ]
  //: joint g6 (B) @(210, 340) /w:[ 2 -1 1 4 ]
  //: joint g7 (A) @(227, 321) /w:[ 2 -1 1 4 ]
  and g5 (.I0(A), .I1(B), .Z(C));   //: @(276,369) /sn:0 /delay:" 4" /w:[ 5 5 0 ]
  //: input g0 (A) @(120,321) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire C;    //: /sn:0 {0}(444,46)(444,100)(358,100)(358,122){1}
wire w2;    //: /sn:0 {0}(188,150)(295,150){1}
wire w5;    //: /sn:0 {0}(186,213)(295,213){1}
wire S;    //: /sn:0 /dp:1 {0}(445,189)(412,189){1}
//: enddecls

  //: switch g4 (w5) @(169,213) /sn:0 /w:[ 0 ] /st:0
  //: switch g3 (w2) @(171,150) /sn:0 /w:[ 0 ] /st:1
  led g2 (.I(C));   //: @(444,39) /sn:0 /w:[ 0 ] /type:0
  led g1 (.I(S));   //: @(452,189) /sn:0 /R:3 /w:[ 0 ] /type:0
  HA g0 (.B(w5), .A(w2), .C(C), .S(S));   //: @(296, 123) /sz:(115, 128) /sn:0 /p:[ Li0>1 Li1>1 To0<1 Ro0<1 ]

endmodule
