//: version "1.8.7"

module CPA16b(S, B, Cin, Cout, A);
//: interface  /sz:(118, 71) /bd:[ Ti0>A[15:0](42/118) Ti1>B[15:0](71/118) Ri0>Cin(34/71) Lo0<Cout(35/71) Bo0<S[15:0](58/118) ]
input [15:0] B;    //: /sn:0 {0}(740,214)(639,214){1}
//: {2}(638,214)(481,214){3}
//: {4}(480,214)(326,214){5}
//: {6}(325,214)(171,214){7}
//: {8}(170,214)(154,214){9}
input [15:0] A;    //: /sn:0 {0}(740,190)(607,190){1}
//: {2}(606,190)(448,190){3}
//: {4}(447,190)(293,190){5}
//: {6}(292,190)(138,190){7}
//: {8}(137,190)(131,190){9}
input Cin;    //: /sn:0 {0}(740,297)(687,297){1}
output Cout;    //: /sn:0 /dp:1 {0}(100,296)(80,296)(80,297)(61,297){1}
output [15:0] S;    //: /sn:0 /dp:1 {0}(722,366)(773,366){1}
wire [3:0] w16;    //: /sn:0 {0}(448,194)(448,262){1}
wire [3:0] w6;    //: /sn:0 {0}(470,337)(470,371)(716,371){1}
wire [3:0] w7;    //: /sn:0 /dp:1 {0}(311,336)(311,361)(716,361){1}
wire [3:0] w25;    //: /sn:0 {0}(639,218)(639,262){1}
wire [3:0] w4;    //: /sn:0 {0}(629,337)(629,381)(716,381){1}
wire [3:0] w3;    //: /sn:0 {0}(326,218)(326,262){1}
wire [3:0] w0;    //: /sn:0 {0}(138,194)(138,261){1}
wire w19;    //: /sn:0 {0}(410,297)(392,297)(392,296)(374,296){1}
wire [3:0] w24;    //: /sn:0 {0}(607,194)(607,202)(606,202)(606,262){1}
wire [3:0] w1;    //: /sn:0 {0}(171,218)(171,261){1}
wire [3:0] w8;    //: /sn:0 /dp:1 {0}(156,336)(156,351)(716,351){1}
wire w27;    //: /sn:0 {0}(568,297)(529,297){1}
wire [3:0] w17;    //: /sn:0 {0}(481,218)(481,262){1}
wire [3:0] w2;    //: /sn:0 {0}(293,194)(293,262){1}
wire w5;    //: /sn:0 {0}(255,296)(219,296){1}
//: enddecls

  tran g8(.Z(w16), .I(A[7:4]));   //: @(448,188) /sn:0 /R:1 /anc:1 /w:[ 0 4 3 ] /ss:1
  CPA g4 (.B(w17), .A(w16), .Cin(w27), .Cout(w19), .S(w6));   //: @(411, 263) /sz:(117, 73) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  CPA g3 (.B(w3), .A(w2), .Cin(w19), .Cout(w5), .S(w7));   //: @(256, 263) /sz:(117, 72) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  concat g16 (.I0(w4), .I1(w6), .I2(w7), .I3(w8), .Z(S));   //: @(721,366) /sn:0 /w:[ 1 1 1 1 0 ] /dr:0
  //: output g17 (S) @(770,366) /sn:0 /w:[ 1 ]
  //: input g2 (B) @(742,214) /sn:0 /R:2 /w:[ 0 ]
  CPA g1 (.B(w1), .A(w0), .Cin(w5), .Cout(Cout), .S(w8));   //: @(101, 262) /sz:(117, 73) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  tran g10(.Z(w0), .I(A[15:12]));   //: @(138,188) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1
  //: input g6 (Cin) @(742,297) /sn:0 /R:2 /w:[ 0 ]
  tran g9(.Z(w24), .I(A[3:0]));   //: @(607,188) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  tran g7(.Z(w2), .I(A[11:8]));   //: @(293,188) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  tran g12(.Z(w17), .I(B[7:4]));   //: @(481,212) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  tran g14(.Z(w1), .I(B[15:12]));   //: @(171,212) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1
  tran g11(.Z(w3), .I(B[11:8]));   //: @(326,212) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  CPA g5 (.B(w25), .A(w24), .Cin(Cin), .Cout(w27), .S(w4));   //: @(569, 263) /sz:(117, 73) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: output g15 (Cout) @(64,297) /sn:0 /R:2 /w:[ 1 ]
  //: input g0 (A) @(742,190) /sn:0 /R:2 /w:[ 0 ]
  tran g13(.Z(w25), .I(B[3:0]));   //: @(639,212) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1

endmodule

module HA(C, S, B, A);
//: interface  /sz:(263, 230) /bd:[ Li0>A(49/230) Li1>B(127/230) To0<C(143/263) Ro0<S(91/230) ]
input B;    //: /sn:0 {0}(122,340)(208,340){1}
//: {2}(212,340)(257,340)(257,326)(265,326){3}
//: {4}(210,342)(210,371)(265,371){5}
input A;    //: /sn:0 {0}(122,321)(225,321){1}
//: {2}(229,321)(265,321){3}
//: {4}(227,323)(227,366)(265,366){5}
output C;    //: /sn:0 /dp:1 {0}(286,369)(380,369){1}
output S;    //: /sn:0 /dp:1 {0}(286,324)(375,324){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(276,324) /sn:0 /delay:" 5" /w:[ 3 3 0 ]
  //: output g3 (C) @(377,369) /sn:0 /w:[ 1 ]
  //: output g2 (S) @(372,324) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(120,340) /sn:0 /w:[ 0 ]
  //: joint g6 (B) @(210, 340) /w:[ 2 -1 1 4 ]
  //: joint g7 (A) @(227, 321) /w:[ 2 -1 1 4 ]
  and g5 (.I0(A), .I1(B), .Z(C));   //: @(276,369) /sn:0 /delay:" 4" /w:[ 5 5 0 ]
  //: input g0 (A) @(120,321) /sn:0 /w:[ 0 ]

endmodule

module CPA(Cin, B, S, A, Cout);
//: interface  /sz:(327, 51) /bd:[ Ti0>A(106/327) Ti1>B(174/327) Ti2>B(174/327) Ti3>A(106/327) Ri0>Cin(24/51) Ri1>Cin(24/51) Lo0<C4(28/51) Lo1<C4(28/51) Bo0<S3(44/327) Bo1<S2(118/327) Bo2<S1(203/327) Bo3<S0(280/327) Bo4<S0(280/327) Bo5<S1(203/327) Bo6<S2(118/327) Bo7<S3(44/327) ]
input [3:0] B;    //: /sn:0 {0}(734,44)(698,44){1}
//: {2}(697,44)(597,44){3}
//: {4}(596,44)(500,44){5}
//: {6}(499,44)(399,44){7}
//: {8}(398,44)(319,44){9}
input [3:0] A;    //: /sn:0 {0}(319,21)(377,21){1}
//: {2}(378,21)(471,21){3}
//: {4}(472,21)(572,21){5}
//: {6}(573,21)(671,21){7}
//: {8}(672,21)(725,21){9}
input Cin;    //: /sn:0 /dp:1 {0}(720,125)(749,125){1}
output Cout;    //: /sn:0 /dp:1 {0}(354,113)(331,113)(331,181){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(256,247)(168,247){1}
wire w6;    //: /sn:0 {0}(500,48)(500,56)(497,56)(497,80){1}
wire A0;    //: /sn:0 {0}(673,86)(673,33)(672,33)(672,25){1}
wire S1;    //: /sn:0 {0}(587,155)(587,242)(262,242){1}
wire w7;    //: /sn:0 {0}(573,25)(573,83){1}
wire w4;    //: /sn:0 {0}(620,122)(650,122){1}
wire A3;    //: /sn:0 {0}(377,77)(377,33)(378,33)(378,25){1}
wire w3;    //: /sn:0 {0}(424,116)(450,116){1}
wire w1;    //: /sn:0 /dp:1 {0}(391,149)(391,262)(262,262){1}
wire w8;    //: /sn:0 {0}(597,48)(597,83){1}
wire w2;    //: /sn:0 {0}(472,25)(472,33)(473,33)(473,80){1}
wire w5;    //: /sn:0 {0}(550,119)(520,119){1}
wire B3;    //: /sn:0 {0}(401,77)(401,56)(399,56)(399,48){1}
wire w9;    //: /sn:0 {0}(687,158)(687,232)(262,232){1}
wire B0;    //: /sn:0 {0}(697,86)(697,56)(698,56)(698,48){1}
wire S2;    //: /sn:0 {0}(487,152)(487,252)(262,252){1}
//: enddecls

  tran g4(.Z(w2), .I(A[2]));   //: @(472,19) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: input g8 (Cin) @(751,125) /sn:0 /R:2 /w:[ 1 ]
  tran g3(.Z(w7), .I(A[1]));   //: @(573,19) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  FA g16 (.B(w6), .A(w2), .Cin(w5), .Cout(w3), .S(S2));   //: @(451, 81) /sz:(68, 70) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<0 ]
  FA g17 (.B(B3), .A(A3), .Cin(w3), .Cout(Cout), .S(w1));   //: @(355, 78) /sz:(68, 70) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<0 Bo0<0 ]
  tran g2(.Z(A0), .I(A[0]));   //: @(672,19) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: input g1 (B) @(317,44) /sn:0 /w:[ 9 ]
  tran g18(.Z(w8), .I(B[1]));   //: @(597,42) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  concat g10 (.I0(w9), .I1(S1), .I2(S2), .I3(w1), .Z(S));   //: @(257,247) /sn:0 /R:2 /w:[ 1 1 1 1 0 ] /dr:0
  tran g6(.Z(B3), .I(B[3]));   //: @(399,42) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  tran g7(.Z(w6), .I(B[2]));   //: @(500,42) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  //: output g9 (S) @(171,247) /sn:0 /R:2 /w:[ 1 ]
  tran g5(.Z(A3), .I(A[3]));   //: @(378,19) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  FA g14 (.B(B0), .A(A0), .Cin(Cin), .Cout(w4), .S(w9));   //: @(651, 87) /sz:(68, 70) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  tran g19(.Z(B0), .I(B[0]));   //: @(698,42) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  //: input g0 (A) @(317,21) /sn:0 /w:[ 0 ]
  FA g15 (.B(w8), .A(w7), .Cin(w4), .Cout(w5), .S(S1));   //: @(551, 84) /sz:(68, 70) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  //: output g13 (Cout) @(331,178) /sn:0 /R:3 /w:[ 1 ]

endmodule

module HS16b(A, Cout, B, S);
//: interface  /sz:(66, 67) /bd:[ Ti0>B[15:0](51/66) Ti1>A[15:0](16/66) Lo0<Cout(35/67) Bo0<S[15:0](33/66) ]
input [15:0] B;    //: /sn:0 /dp:1 {0}(524,257)(524,242){1}
supply1 w0;    //: /sn:0 {0}(620,351)(620,336)(572,336){1}
input [15:0] A;    //: /sn:0 {0}(495,249)(495,301){1}
output Cout;    //: /sn:0 /dp:1 {0}(452,337)(407,337){1}
output [15:0] S;    //: /sn:0 /dp:1 {0}(511,374)(511,405)(464,405){1}
wire [15:0] w3;    //: /sn:0 /dp:1 {0}(524,273)(524,301){1}
//: enddecls

  //: input g4 (A) @(495,247) /sn:0 /R:3 /w:[ 0 ]
  //: output g17 (Cout) @(410,337) /sn:0 /R:2 /w:[ 1 ]
  //: supply1 g2 (w0) @(609,351) /sn:0 /R:2 /w:[ 0 ]
  not g1 (.I(B), .Z(w3));   //: @(524,263) /sn:0 /R:3 /w:[ 0 0 ]
  //: input g5 (B) @(524,240) /sn:0 /R:3 /w:[ 1 ]
  CPA16b g0 (.A(A), .B(w3), .Cin(w0), .Cout(Cout), .S(S));   //: @(453, 302) /sz:(118, 71) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: output g15 (S) @(467,405) /sn:0 /R:2 /w:[ 1 ]

endmodule

module main;    //: root_module
wire [15:0] B;    //: /sn:0 {0}(234,170)(234,139)(312,139)(312,116){1}
wire [15:0] A;    //: /sn:0 {0}(199,170)(199,140)(121,140)(121,118){1}
wire Cout;    //: /sn:0 {0}(182,206)(99,206)(99,404){1}
wire [15:0] S;    //: /sn:0 /dp:3 {0}(349,398)(349,347)(218,347){1}
//: {2}(216,345)(216,239){3}
//: {4}(216,349)(216,390){5}
//: enddecls

  led g4 (.I(S));   //: @(349,405) /sn:0 /R:2 /w:[ 0 ] /type:1
  led g3 (.I(S));   //: @(216,397) /sn:0 /R:2 /w:[ 5 ] /type:2
  //: dip g2 (B) @(312,106) /sn:0 /w:[ 1 ] /st:22
  //: dip g1 (A) @(121,108) /sn:0 /w:[ 1 ] /st:26
  led g6 (.I(Cout));   //: @(99,411) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: joint g5 (S) @(216, 347) /w:[ 1 2 -1 4 ]
  HS16b g0 (.B(B), .A(A), .Cout(Cout), .S(S));   //: @(183, 171) /sz:(66, 67) /sn:0 /p:[ Ti0>0 Ti1>0 Lo0<0 Bo0<3 ]

endmodule

module FA(Cout, S, Cin, B, A);
//: interface  /sz:(169, 168) /bd:[ Li0>A(43/168) Li1>B(84/168) Li2>Cin(126/168) To0<Cout(98/169) Ro0<S(83/168) ]
input B;    //: /sn:0 {0}(125,198)(216,198){1}
input A;    //: /sn:0 {0}(125,181)(216,181){1}
input Cin;    //: /sn:0 {0}(132,107)(277,107){1}
output Cout;    //: /sn:0 /dp:1 {0}(391,153)(419,153){1}
output S;    //: /sn:0 {0}(299,98)(299,67)(317,67){1}
wire w1;    //: /sn:0 {0}(239,175)(239,155)(370,155){1}
wire w8;    //: /sn:0 {0}(259,199)(269,199)(269,121)(277,121){1}
wire w5;    //: /sn:0 {0}(319,114)(360,114)(360,150)(370,150){1}
//: enddecls

  //: output g4 (Cout) @(416,153) /sn:0 /w:[ 1 ]
  //: output g3 (S) @(314,67) /sn:0 /w:[ 1 ]
  //: input g2 (Cin) @(130,107) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(123,198) /sn:0 /w:[ 0 ]
  HA g6 (.B(w8), .A(Cin), .S(S), .C(w5));   //: @(278, 99) /sz:(40, 40) /sn:0 /p:[ Li0>1 Li1>1 To0<0 Ro0<0 ]
  or g9 (.I0(w5), .I1(w1), .Z(Cout));   //: @(381,153) /sn:0 /delay:" 4" /w:[ 1 1 0 ]
  HA g5 (.B(B), .A(A), .C(w1), .S(w8));   //: @(217, 176) /sz:(41, 40) /sn:0 /p:[ Li0>1 Li1>1 To0<0 Ro0<0 ]
  //: input g0 (A) @(123,181) /sn:0 /w:[ 0 ]

endmodule
