//: version "1.8.7"

module HA(C, S, B, A);
//: interface  /sz:(78, 65) /bd:[ Li0>A(13/65) Li1>B(35/65) To0<C(42/78) Ro0<S(25/65) ]
input B;    //: /sn:0 {0}(122,340)(208,340){1}
//: {2}(212,340)(257,340)(257,326)(265,326){3}
//: {4}(210,342)(210,371)(265,371){5}
input A;    //: /sn:0 {0}(122,321)(225,321){1}
//: {2}(229,321)(265,321){3}
//: {4}(227,323)(227,366)(265,366){5}
output C;    //: /sn:0 /dp:1 {0}(286,369)(380,369){1}
output S;    //: /sn:0 /dp:1 {0}(286,324)(375,324){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(276,324) /sn:0 /delay:" 5" /w:[ 3 3 0 ]
  //: output g3 (C) @(377,369) /sn:0 /w:[ 1 ]
  //: output g2 (S) @(372,324) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(120,340) /sn:0 /w:[ 0 ]
  //: joint g6 (B) @(210, 340) /w:[ 2 -1 1 4 ]
  //: joint g7 (A) @(227, 321) /w:[ 2 -1 1 4 ]
  and g5 (.I0(A), .I1(B), .Z(C));   //: @(276,369) /sn:0 /delay:" 4" /w:[ 5 5 0 ]
  //: input g0 (A) @(120,321) /sn:0 /w:[ 0 ]

endmodule

module RCA2b(S, B, A);
//: interface  /sz:(40, 40) /bd:[ ]
input [1:0] B;    //: /sn:0 {0}(123,112)(195,112){1}
//: {2}(196,112)(300,112){3}
//: {4}(301,112)(322,112){5}
//: {6}(323,112)(506,112){7}
//: {8}(507,112)(535,112){9}
input [1:0] A;    //: /sn:0 {0}(123,89)(190,89){1}
//: {2}(191,89)(295,89){3}
//: {4}(296,89)(317,89){5}
//: {6}(318,89)(501,89){7}
//: {8}(502,89)(534,89){9}
output [3:0] S;    //: /sn:0 /dp:1 {0}(121,346)(68,346){1}
wire w13;    //: /sn:0 {0}(504,175)(504,331)(127,331){1}
wire w6;    //: /sn:0 {0}(296,93)(296,154){1}
wire w7;    //: /sn:0 {0}(308,283)(308,341)(127,341){1}
wire C0;    //: /sn:0 /dp:1 {0}(187,282)(187,361)(127,361){1}
wire w4;    //: /sn:0 {0}(320,203)(320,175){1}
wire w0;    //: /sn:0 /dp:1 {0}(191,93)(191,150){1}
wire w3;    //: /sn:0 {0}(203,282)(203,351)(127,351){1}
wire w12;    //: /sn:0 {0}(502,93)(502,154){1}
wire w10;    //: /sn:0 {0}(318,93)(318,154){1}
wire w1;    //: /sn:0 {0}(301,116)(301,154){1}
wire w8;    //: /sn:0 {0}(193,171)(193,202){1}
wire w11;    //: /sn:0 {0}(507,116)(507,154){1}
wire w2;    //: /sn:0 {0}(196,116)(196,150){1}
wire C;    //: /sn:0 /dp:1 {0}(268,240)(252,240)(252,187)(215,187)(215,202){1}
wire w5;    //: /sn:0 {0}(298,203)(298,175){1}
wire w9;    //: /sn:0 {0}(323,116)(323,154){1}
//: enddecls

  tran g8(.Z(w6), .I(A[0]));   //: @(296,87) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  tran g4(.Z(w0), .I(A[1]));   //: @(191,87) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  HA g3 (.B(w5), .A(w4), .C(C), .S(w7));   //: @(269, 204) /sz:(65, 78) /sn:0 /p:[ Ti0>0 Ti1>0 Lo0<0 Bo0<0 ]
  //: output g16 (S) @(71,346) /sn:0 /R:2 /w:[ 1 ]
  concat g17 (.I0(w13), .I1(w7), .I2(w3), .I3(C0), .Z(S));   //: @(122,346) /sn:0 /R:2 /w:[ 1 1 1 1 0 ] /dr:0
  HA g2 (.B(w8), .A(C), .C(C0), .S(w3));   //: @(164, 203) /sz:(65, 78) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 Bo1<0 ]
  //: input g1 (B) @(121,112) /sn:0 /w:[ 0 ]
  and g10 (.I0(w9), .I1(w10), .Z(w4));   //: @(320,165) /sn:0 /R:3 /delay:" 4" /w:[ 1 1 1 ]
  tran g6(.Z(w2), .I(B[1]));   //: @(196,110) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g9(.Z(w1), .I(B[1]));   //: @(301,110) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  and g7 (.I0(w1), .I1(w6), .Z(w5));   //: @(298,165) /sn:0 /R:3 /delay:" 4" /w:[ 1 1 1 ]
  tran g12(.Z(w9), .I(B[0]));   //: @(323,110) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  tran g14(.Z(w12), .I(A[0]));   //: @(502,87) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g11(.Z(w10), .I(A[1]));   //: @(318,87) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  and g5 (.I0(w2), .I1(w0), .Z(w8));   //: @(193,161) /sn:0 /R:3 /delay:" 4" /w:[ 1 1 0 ]
  tran g15(.Z(w11), .I(B[0]));   //: @(507,110) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  //: input g0 (A) @(121,89) /sn:0 /w:[ 0 ]
  and g13 (.I0(w11), .I1(w12), .Z(w13));   //: @(504,165) /sn:0 /R:3 /delay:" 4" /w:[ 1 1 0 ]

endmodule

module main;    //: root_module
wire [1:0] B;    //: /sn:0 {0}(155,160)(155,202)(237,202){1}
wire [1:0] A;    //: /sn:0 /dp:1 {0}(203,130)(203,167)(237,167){1}
wire [3:0] S;    //: /sn:0 /dp:1 {0}(294,265)(294,241){1}
//: enddecls

  led g3 (.I(S));   //: @(294,272) /sn:0 /R:2 /w:[ 0 ] /type:3
  //: dip g2 (B) @(155,150) /sn:0 /w:[ 0 ] /st:3
  //: dip g1 (A) @(203,120) /sn:0 /w:[ 0 ] /st:3
  RCA2b g0 (.B(B), .A(A), .S(S));   //: @(238, 138) /sz:(111, 102) /sn:0 /p:[ Li0>1 Li1>1 Bo0<1 ]

endmodule
